`include "svlogger.sv"

`define ENABLE_DUMPVARS
`define DEFAULT_LOG_LEVEL  `SVL_VERBOSE_INFO
